//ALU testbench, just test using CLA through ALU for now
`timescale 1ns/100ps
module ALU_tb;

	reg [31:0] A, B, op_sel;
	wire [31:0] Zhi, Zlo;
	//wire[63:0] Z;

	ALU alu_inst(A, B, op_sel, Zhi, Zlo);

	initial begin
		A <= 32'd0;
		B <= 32'd0;
		op_sel <= 32'd0;
		//Test Addition (works)
		#10	A <= 32'd8960;
				B <= 32'd6500;
				op_sel <= 32'b00011000000000000000000000000000;
		//Test subtraction (works)
		#10 	A <= 32'd80000;
				B <= 32'd10000000;
				op_sel <= 32'b00100000000000000000000000000000;
		//test Multiplicaton 
		#10 	A <= 32'd960;
				B <= 32'd60;
				op_sel <= 32'b01111000000000000000000000000000;
		//Test division 
		#10	A <= 32'd8;
				B <= 32'd3;
				op_sel <= 32'b10000000000000000000000000000000;
		//Test SHR (works)
		#10	B <= 32'b00000000000000000000000000000010;
				op_sel <= 32'b00111000000000000000000000000000;
		//Test SHRA (works)
		#10	B <= 32'b10000000000000000000000000000000;
				op_sel <= 32'b01000000000000000000000000000000;
		//Test SHL (works)
		#10	B <= 32'b10000000000000000000000000000000;
				op_sel <= 32'b01001000000000000000000000000000;
		//Test ROR (works)
		#10	B <= 32'b00000000000000000000000000000001;
				op_sel <= 32'b01010000000000000000000000000000;
		//Test ROL  (works)
		#10	B <= 32'b10000000000000000000000000000000;
				op_sel <= 32'b01011000000000000000000000000000;
		//Test AND (works, bitwise)
		#10 	A <= 32'b00000000111100000000000000000000;
				B <= 32'b00000000111110000000000000000000;
				op_sel <= 32'b00101000000000000000000000000000;
		//Test OR (works, bitwise)
		#10	A <= 32'b10101010101010101010101010101010;
				B <= 32'b01010101010101010101010101010101;
				op_sel <= 32'b00110000000000000000000000000000;
		//Test Negation (works)
		#10	B <= 32'b00000000111111110000000011111111;
				op_sel <= 32'b10001000000000000000000000000000;
		//Test NOT (works)
		#10	B <= 32'b11111111111111111111111111111111;
				op_sel <= 32'b10010000000000000000000000000000;
		
		#10 	op_sel <= 32'b00000000000000000000000000000000;
		
		#10	B <= 32'b00000000000000000000000000000000;
				op_sel <= 32'b10010000000000000000000000000000;
		end
endmodule