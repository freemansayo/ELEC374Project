//acts as Top-level design object, holds the control unit and datapath modules, facilitates communication between the two.
module MiniSRC();
	
	control_unit CU_inst();
	
	Datapath DP_inst();
	
endmodule 